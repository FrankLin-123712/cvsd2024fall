// list all paths to your design files
`include "../01_RTL/core.v"
`include "../01_RTL/system_controller.v"
`include "../01_RTL/sram_4banks.v"
`include "../01_RTL/sram_bank_controller.v"
`include "../01_RTL/conv_engine.v"
`include "../01_RTL/sobel_nms_engine.v"
`include "../01_RTL/median_filter_engine.v"
`include "../01_RTL/four2oneMux.v"