`include "../01_RTL/define.v"
`include "../01_RTL/utils.v"
`include "../01_RTL/ed25519.v"
