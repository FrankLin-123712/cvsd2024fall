package dat_0;
integer pat_num = 0;
reg [767:0] input_data  = 768'h259f4329e6f4590b9a164106cf6a659eb4862b21fb97d43588561712e8e5216a0fa4d2a95dafe3275eaf3ba907dbb1da819aba3927450d7399a270ce660d2fae2f0fe2678dedf6671e055f1a557233b324f44fb8be4afe607e5541eb11b0bea2;
reg [767:0] golden_data = 768'h2f8a66a8da71da5f8c006b1aa2fd5320e6dab0b39ff360b34fe039289869012545a22939c0fc3f79f416185ad1e5404ad7266f50b66617b28733045dbbf700a252310c49eea9ed11b646027438b6ae9e7e7885841a35ed71e541e372bdd37189;
endpackage

package dat_1;
integer pat_num = 1;
reg [767:0] input_data  = 768'h17e0aa3c03983ca8ea7e9d498c778ea6eb2083e6ce164dba0ff18e0242af9fc32e2c9fbf00b87ab7cde15119d1c5b09aa9743b5c6fb96ec59dbf2f30209b133c116943db82ba4a31f240994b14a091fb55cc6edd19658a06d5f4c5805730c232;
reg [767:0] golden_data = 768'h7074238c34bf23a70a4eb431e085dd6e83f54385c101e15b04a02078e25e169c573b99fd279b58c07c642837f47d5ffe2e94f81a92d111af2f134f44a1d24d1c3966bdd9ab22ad41aa04ada33003ad2511a5920b3e9c6f395f952374ca68549e;
endpackage

package dat_2;
integer pat_num = 2;
reg [767:0] input_data  = 768'h1759edc372ae22448b0163c1cd9d2b7d247a8333f7b0b7d2cda8056c3d15eef75b90ea17eaf962ef96588677a54b09c016ad982c842efa107c078796f88449a86a210d43f514ec3c7a8e677567ad835b5c2e4bc5dd3480e135708e41b42c0ac6;
reg [767:0] golden_data = 768'h63356304fcc5389ca4b720b26a05d63d7581446982ef76b69da9a536727f3a16360dda0bf1f554083eaa052949519b91d5b0bab0fc8ac857cde46c7d2b13e671785890ce4f71ecb7ff5d8ce5458bd3e0e8edb7718af4bf0ee2142fd45eedfe20;
endpackage