// list all paths to your design files
`include "../01_RTL/IOTDF.v"
`include "../01_RTL/SystemController.v"
`include "../01_RTL/DataLoader.v"
`include "../01_RTL/EnDecryptCrcgen.v"
`include "../01_RTL/Comparator.v"