package test_patterns_pkg;
    typedef struct packed {
        reg [767:0] input_data;
        reg [511:0] golden_data;
    } pattern_t;

    parameter NUM_PATTERNS = 100;
    const pattern_t test_patterns [NUM_PATTERNS-1:0] = '{
        '{768'h099c1716690dae84f20d267415c01fc0b2994f2dc8a7e19eaa136241fd7583257dd22e224f3ba68e8a2b2eb1673772d8aa1a791122c2f3b09be44dea333169c01bbab60da5bfb99594908b631a031effef8005340706003690bf8c4ca0e26f1a, 512'h5643ba63f2518c809870a630ee3ee91d66d20536c5795d714dc416394ed2dc40513fe9ef07a2e7537f6931d1c562b8dfccbd7d191d30ed55f94492a7b3665d34},
        '{768'h494f6bf2e4d4ae140988303d9cf4914f602c3d65026ab837abf7d55b0bcc80e015107d64851b646122bea321345d74d75d243984905d1e46ec0c866a667556bc1ecaae4512dc15cc91781af297ae9496c2158be4225d17ad53f9327d714c7c6e, 512'h14ea66c12ea72baae24f2ee47c7d6bcaeebcddcbfc962837def2eff3f7a66c60391d88cb9c64a2145dc6440408424ab58e325f6e3dbff780f7da95f9656b0ec2},
        '{768'h58cb3a607d0abc20a9999c2852b498efe3aab86fbc2eeacee24eeb4b4af0131370deaf169ceddb0195056ccd30097201bb8dbd756b047a98cb927e871699c0db782d08586b924557d14610e049ee0ddbcff6b0bb920602446c054888f72d4c8f, 512'h6e114f9c80b118c9f0a906b1ae069f4f2aa2adc8dc2c59cfb65b02711a1781c8270a5d78b835d3a3cf8614755c25d6b7ce92a052d382e7f1f94f5362a8fb60c2},
        '{768'h42770e34250193ff8095d1096005f425eade8660bc81aa833670d33f946091df277ab780086acf261b0fa1deced1379945f10c69ddfb2f14971a77171886a8456cd1305521b6e2a056bd76de9acbaa408b031412f248a8e6d5909a00fe44d5ef, 512'h21714f36b9eb0801e6ee847d087562ce552e58ee8a17b93910143d517ba1d6080ad1cd162ad150611ca71efec0b6998aa5c78e6e24ea683332feede0fda7112e},
        '{768'h45ab0c1fb9beefe9aa8372a31d6427f1f7a62f7ca07e3845ad5c81bee692a87e2a653e5a863b3070e07dfc577b18fc32c06d2b63adaefe4ee49f1afe86d96e3f668b77d0420fe1cd7e77e5940e06c02f5cd7cd23990fad5e995c031402e80063, 512'h0cf337e45c679c659b581724a3821e7731a113ba89a257d539961009a0c574b228caba2f8892cbdd6850b9abdfac1cc33b606739bb09cc19f3a00a407e0f82aa},
        '{768'h5ca4639fd0a82ba2a2722078db5befdf7f55f5ff52290c512e4cb5e816763e6b04bdd767e735de8a791dd63e5e68d482c1472232915e6c7c976dd11bcbd2c1846e5e304bb0519314b18430b13c4a53e3a9676789e6bd679b6cfbec798157e758, 512'h0dc210bbe4ee3c64cbc2be84034486bf1a6ab36f762e47da05ddc17e09af9c524bd0389d52cfb51c48d7bd3768c4208e02b60e40514b6099f65679feb727d7be},
        '{768'h3c1f9f1f609cd0630d2c45be7af9bf7331b41b907453247b2e0b435b6d57fbc81a2ae727b73a8ffb1852de94aa85c33088cf24998c8eee17dc9a22c71a51f4186d450563965913bdda203f4fb0ac4226b81b224475f5609b8bfbee54e9f7ce22, 512'h69d4d1ac991d8263a25578dbc8795ed1dd58e6aa8c887af9e935acb7930a912a4bdb119a89b2938bc52f55e799bfdaf686dfcc7b550fac7432f773fe63f9983e},
        '{768'h203717a2e2149d231dcdfe44cbed142b9bbeb17fac761e84a4f99aaef7ac0d1c4f6ee4aa6533f881ff94467bac137dcba284dc20ca7aa2a52b22b791631f91a606ec53ed2c93265f0e2282736836cf7db60acf708bedfa3c6feb03a307c6eb4a, 512'h1888e81e5e2029bb89645b2e168ac71a95a1bfb5abd54f3a01f7efd173be65f214d180839937bfda6116d85337e277406f2abda9b1579838dd88285b8ad46be0},
        '{768'h63464405410ae9da7781b3f39a74797a6e52d39b024ffac30d7b383615d5fffb2951d5ebcb711614c957dc6d7bfc37173ed8e725af0416acd7a686ce8a605e786384d8864cceef180c8cd3fda3a20afd930b657a43fd5f9504188719ee8d0f4d, 512'h4e0d726210441feea2901ea9bef344679419bc7189be83fd66b52afd9a1bd5b834601b71f1af1ab7ca7ee13cdd4ff18faf97332be87a938cbbfd02021214d174},
        '{768'h542e35b68a8ab356fe335aaa577f08d3dcaaa97716bb8bde55f72093a99284163801fcb95461735aadedcf8d019765701768f1eddd85bef5c61d41f814b4a0980f6182ae94ba2b01ad5613e3f827a55e1317661ef89cba33e0b8b599f8873a09, 512'h4c39e436f81288d605e8f74484cca8c338167cfbc20ae3fa34c9d9408957abf65ce2b1a39e4a7351b1e17f3056164f94e4a22c1ac572c1067a2ea35896288646},
        '{768'h3d12115dfd8bdf875a890470996d4d0ed4b93879034de809b8117dc3faecaeee1735bf49b1baba82c49ba482c8338db4d91f0dbe8ca40d9944bd758a3c40be7526da17c3ded1d88bb8e3e0f25349754923d86846cdcf71c043e1265ff1aa9f96, 512'h1afcd5b033df2163cbbda454be39ae53c2accb21a4dda2d976e409dc1c90e4fe002c7ba18a5b54cbaa387cace8f7c828e1e138531450429e4d58a977c183b20c},
        '{768'h04e0c08fa5ea5e1b3b30ab78c6ef0f886d665eaa3c38ea160495f667f5d4f17a5aae0834016ee03b4e2d5a4751043c63581b6b6a7596d9a81dd45b4510bca4670b3287fadeb4d0191739664ea37a8661707ea104eccd8118ebd83a7f085bbb87, 512'h27be6c3031bd7be5b76210d3599058e7850f4a846d861cf8428fdda72a057efa5406aa1d3a9172ee4c53462d41a8f765d4357dee46d2e4b63a1e5ed4c1794f24},
        '{768'h361e326c95b89e33236dc4944a24c9617a67243b90cb9e6b58c7b203265ab2d46231a7f4d18024237e579d9581c3eaa0f412d0771a02453a022216d80aa9f4040acfb37cbafdb4bc9ad19dd5a8fd53394743e54c61e0501958289c6b1b35f71b, 512'h2fe6f720d997520363cbcfaca67d7fba676db44fccf96cf44ebfca020147bc64128c8fde643a48c876af9381962bced2e1e78845c2963dcf472abf16e5cc417c},
        '{768'h2cae122a66ef4554bd26535eac740917267ef7469370d39d44bea6fa12d44b8a7ed1d53c640862462a7f5e299dd365214096b213e6cc6b74bd724369ca630c730ccd3f9b3a1f5ca98d96eaa257f577ddc6efaa523fb337293dde29b2abdc7bb5, 512'h0cb71670582172784e7759f1eb3814d9944cbe087fbcb196769914e256e254ca0bb83133ac61856f0f2aec7cbb3765e0a1c57c54199144073085da024e93edf2},
        '{768'h763e773f2e0c2f528227544b8d9ac17cc3e7ccf8d405daeb7db673c762e836fd70f60c6c86f81a2bedb5bbf0ee1e47e53ea291671ae0111e9c924d5981bbd6ee6959e53e532c008b9e03e24d0ade5577700f1600143ae36f43ec798e47e197f7, 512'h18b4df4c694f2888391c4e6715e40904fa539ef669dc52864d457c097e7857e057307a5e92637e411df5cda6829c02380663d21e2a0e637efa8c5adbe51eae08},
        '{768'h5259669f572b53d555fa8e9c6370d1019cdf9bfb2c3a03407d4168417dba0aef67f2078a50a64c3a2fa27ceab48108dd14aeac45b0fe5f70f15e3176f4bbc07d6329c7b19fa56c8da55be7c1669197361898865a1b29764230d5803f457020fe, 512'h092e3df3597c1deabc67274e1fd10ba4d5ab84014949a7d74800eea20a560f3e6e1a7bcc33dd34001ec779dcd5f7d8bb1c1f8376fd4709a5ac9ba90ebfdabf88},
        '{768'h201929113eb2b7c5da9b1084ef2a88258c3a2bbf8365e0afdc8766b4a6471a9053226254030dfc34901d39896594e44a15e511c89990bda65b8db5b0f4ef80dd4a5be027235d46551831a59973a198ec577a45576017fa017101a860f30a1405, 512'h4d0e77226fa8049200ce834f028f37813ae1f59fa00f8609cba3621e45f5c9a06fdda22d74ee360d5c040b931f6dc31d0247eb9d72f66d01570c5ce84cb25344},
        '{768'h46df1f9eeff09e8f2ae2cc58c4419c4a5397a7003414ab5f932b662cd640ec2464643557ba5709502657a91c4e6659d312f7c018170d1882da9ad1aca8f41f60125f1a29ffdc2c356f1e230b4d0de574806936b77cb2daa2a1f4150a259a7fc3, 512'h27eedf69d20500383fa8b89cc686e8be1aaaf691f198cab221cf1df3dd99d50428ac15c6abf78af58536eb2fe11bd572d9a0326b53e34f5aa905315ffdb404c6},
        '{768'h3c44c17c83f385d99d5d40d9b8fbbc5ffe426bb4c8f457b722a1980acb5a00782165f308bf0c09651d45f6e68f611b2676fc103ce830e783cde6b02ec32f9f757def13d7bd297cc29b9c862d52ef90ee5e51701b4c548d2c7226a470e466d4b6, 512'h73f804b568fbfae33bba49c7b7148baa66f8459f506390cb288957bc8b9b457e0cbaa95cef35b042f19fe8941b0ee0811baf9517a1d7c7ad4251c3f2e99c1a7e},
        '{768'h38221fbe4b0f8fc85dff39c49f639568429d28b9a451d27d993a65e1711c1fac19ecc79d321c0cc0d13c1c5a21a77095a546b05a3036ad08622d2f291c35e7760577371ce022b1799859bd89a0eb4e50cf853b8ffdc78d23b27e17ccf421857b, 512'h1060ad7aa77aa44fe9b4bb1a52c8f0e9ee7074d8dbb08d8bc17a2fcb58b449b2142af1369141ac457373b2b59f9b77a0977b7416ba5e26e0508f96505e9e66f0},
        '{768'h479adcf5c895e46e7a56c54fce0c806b003086522d276b4dc657bc1e3978a75266b4bd82c0d04baa86a71418d6c82559d5f84a7aaeedca2e4dce96d6d41605d51b0c1ebea3edf95af9ab5257dea909270869ec63c8f914a1858a951ea23bcbf2, 512'h6da395b4bc82d3466c9d9d1e021e7614d5bdcf61223f5fd85fa30edfbab1e1ba0f9a0f831540ab7ea61382d71585c5e581ad6baa5ed4965bbbf761ef439d6344},
        '{768'h1f290f09e14a894d120b9f1706687fb666bf56bf0e52b542accfec3c7a8f49f35a061fb81906c932fe9d1f907dd2b2488c6bec7f3f3b417ad275dc67cb51761268ca0a2d600873b0e5de08836c73f77e7473cfb68b601c0d603e90f068cecb90, 512'h7ce5d202cc36b5f86b402e1f580b49e560de3dd91f9e333375fb40452b07cade41c891b0d7fe92bf25befb5064b00faa06bf2ff317836d7a97ef5de4b27e5c84},
        '{768'h436289697de9022af287129bc2f2915053c7ac3f7d18244d2d75e6855835671a29509b0865d968269360dd3401745e2eb0d24f6233a0a4fbe1fcb806d64d33ab0083ff5f7c3eb427c17ccc0872bf56fbcb8e79c7b224208f79bf3ca874644a4e, 512'h27a2fb36f2bc2dbc321dd2b6f7fd88da0794f09981f86d8045a37d30a883996c5324f02418b2a107896eda0de7ed275218c94120f76b3149d8d567b5d6ee1efc},
        '{768'h5e24681c74c6f5792701e55608e1a7b5cf7a76337fa674907a789301dae636786709ff744d1f9e53401d754752dd4349ad1d0436333309e1d0e0ad7248af50322f7a8b2375d32c6ca27eea4a5c294ad5b92a8a633a1751f37c5b59ecc369fba9, 512'h7e8979743ccb79d63b601635ebe90560ec3161c0c2f6c91736b99f984ba032ba773f2f31bd33bf9c89d45e84d8baacd6b90acfd6618b00447bdb6a05911557c4},
        '{768'h6d104e595e1075bec9d5784674a52911a4ecfcc03bb4eb344e25d2443fca021b1988ce840bcb795978f189c4b01753665d4d033ba1587b649d81f3c726025305766480299c011573f5323b4a61c44254af64ccc06c553c1975efac2dd364f8b4, 512'h6aa168302d680658666fc55313066076971ead39810a47ea8f3f298543676b964c13fb2c92ca7f6da4318d25dda13fce7a2690c96aedad28e5102da9bed43840},
        '{768'h0a7ed65d7312391c21a9d5fcd66be6f203b1e11256afb025027cf9e086fe7eb6401cb540cfc2b2ac0f1c6227bc31a161af885805f8822328c893c97c7d629f531b72eb4bda9d1d384f96280a0dbae8c1e1b659f7e80ba1789a2df4fd4bc9ff1f, 512'h7ae39380e1633e63724b7b9c364518b592d799ed522221e82a7a1e36958b663a3d1d6b225ba689dc39dbb536d2f198d1d0dd9e660d0ebe551d65902b1a57539c},
        '{768'h41c1091998224564fb389b45a7f5b759fd2bae1191181bc1a27ce9e7b41fe0a34489f7438ae8760dbcde2a10579410a3fbeb82b24ef8cefbbfbbc02bd108653871c75546830a4a48cea6204372488e083e0541d581813d4628bcafdccdca719c, 512'h1be04bfbcec9fb0b0b7116fa08b20cea4fd3da4604ea2dd6c34de5c9b68f16d23227ae19d119080bf5093beb24e748d72daf91c02a6d5e73f1f571a878d2a5f4},
        '{768'h77edf92b4ce14600ede4edee6d0568aa00f54404695709d5f6afe310cd41c33a6521510b7043fd77e4a16d28831a919ba05085b2b39b74267f35154135d11e6724cea083ed923752a357fae285939168ce954a0deaec32a9a9ee6451abed02e8, 512'h57c5de46af894d8e5951229ba71856278831264300988110e0cb1bfe88610faa4b579457db440251fee2c7183bc729f4658aeb105638e81e78aec6856eb8cd5e},
        '{768'h52d6731dbc6f01f19c72e9c2d05fc8c00e2bac4b0a082986aa06ffbf32eb062b685c39aa10259bbbcf285a29df56e6d84386cc14045f3ab2b262cc8f25a759642e87be33c486e15fd5af594858b4936248a9d461bd943d315c0dfbe1d2d1e82e, 512'h61b3a3d760453a4c1905d340787f9744d8652465374613651958f0eb9331ff2a37e6021f561bff7c517b352eacc0002ac6de9d2ae8b1ab13c4bfb1af840244ca},
        '{768'h6b2a9ce37912017897ffbdad568846becd7b981263cf6b1bbc8cb07220ce65fe05ef249997a2de73a189f5d681e79f70dc7cdff02f11dae1aefb916b99c0a3ef5941daaed9108b8e94c3210f9a57088931489eccb504b83d80c799512ba0d4e9, 512'h401b73a2172a4acd7241fef1247c1c53411a7d70748b2b1062bde1e7cb60b1aa7e76b1bd045e2e939d42d6df7c05ad7695cd8576aff600b965378241990d6c86},
        '{768'h0814715b8283fb6661720f9eff2a29c4198c0456a462ae0a8fdff72591a71b0b1d185603b376c8f58786a8c4eced506ac1e39ccbd6cd90927db39880e11e3a3043a3822824f66a3642f44b130104c342aa95e47e18f88d6ef22ef63618b365da, 512'h363f43149379ee82101302a757642764f6683a836f71812b41d8383c98f8d7f07205d8e84aeec0700faed5f1b81c0ff990593effd282b7abc5cf6cc8aaea23a0},
        '{768'h011f522f9fbf610562d39fd380b07263dec4294a9e23335b2bf1e6c5894b0e5b6a3b22e7eba0c65b5e14c9b4480dd51d62782aba4f8ca2b3b7be91a5c594693e620cfa894043c895db0cc9251c9774de7d54fa7ff98f44dc0581339429f78d23, 512'h0d2c05fd48b6708710def50d8d56fb574806074d66fc9c95da72ebce26a73bf82020f84498f7523ba6f288b870ce172cc71ebbe5fd7080af1c1d08e775415474},
        '{768'h27f2f2b0781525407693ae6264c69629d4fd7b5c7f96d8ae8bf18aa1fdede45752036635141d6c5d0cc0c4647bceda6113866ac82e2a4e2dfe9bfff2f03d7c86684d097109ca4341653f88e7b4306eb8260d44d5e80ceee8adfdf5490c8bcabc, 512'h32275890f70b8d0cf9deb7be5e2c9f7f52fb1e7e3f256e6c40f81d04de63389615e21a685debd18c807c5ac64184832cae13ba8be8c612a67493af307f095162},
        '{768'h7f752c76da58e54f4000528c13d8047aa1fac106803c6adac2b1018943569d0a3b714a1dbc15c94886cc2d73f7c1f7645e4a5d7f02748f87b7c150ec88edc6a82814d81ea6ce889fe78d7d17ddb01d3fff0c541fc080622643c4ec947e656d51, 512'h1c5898607149fcad1b819a243fce5680169bffd1c2b7be88f5b50f51ffe25e0a3a25b94f1a201f944e74fa1781f1df0b3f1fc79a6695cd8e330f585a71382a44},
        '{768'h348653c1fc88d751f114088d331ad631be4918c0e14eb42124bf02d92bf6b7067fc2bcf63b787193888ef620ffab25f0eb5b17f57fe79b81fcec4a3764b00bfb26c9b051d86497a6d222eec5cba2eb226f2254a6d8f21b08cf0a08cf26122c17, 512'h08b998d1fc91e2f03d272a67ebaca39ee5856a6886588247217fc652637d479c16ec4df6b373971fce817ae8c81c2d8f1442838087a24ab08760b3f8563fbc44},
        '{768'h1cfe168d5b3d5f0e7ee76ddf4691ee1ae0db512152fd04ec3648804996bf7892264f9fe86549f5419f9e9e7885eafcf183ac1759c9d782ffcc8b2918806a0b087c9ad7af629e61973cee3b41a15a948676f57e3dbfe0eea723c21b3f6d9167ee, 512'h6f883f6bb0af1c5842841b502a2169598dd2fab3137a3b4d9d262fb230a0bb26103e4fa87679265941d5af204edb23f48125364d30f0a2bf68da1f460c2f64aa},
        '{768'h30cc60171c5444f719ec69aa982b783de6271c43376a3ee26381a4731a99a16000e2b46b7447ff9e79ce5c94fa39b3d723230251c75882b3f23f7c6780e74c277e4adc4395b7d65e4b040d49cee8fdb867813d0ebc4ba27d1666ba3ba7b21e1e, 512'h054cf3e0988a724fe7fb025da0a1fdb48a97a8c006639b05b787a7a03630c3f01e6a0829a8751cd091f7de70495c8d369a2cea7a8e5db6c62be70c6eef1da4d4},
        '{768'h450e2945defd2370d3f7d3c330c569c51e712f37c2481a1f48a4bd0326cdb8001976433df1fd7d03261c85ca573d71086c1fc81746c1eb9985cddc61b90e7e1b2effb8668112cf0fd3bafeefb9b7068fc423c4074a71025de17be0528e21f3fb, 512'h2a64f7a41df78d95f10ffeb8f43652350354cbba81d14a1c218b3a472fdf743a781efc41ca757fc863e177090e4a38d7159846c440be2ec20bfcb6e668bf76c0},
        '{768'h4fdaec2be4008005ce205ad6dc0e399bf8c32ddf3107d6c922f57caea445ac623476dd6707602320c5f9e28d05a4a8ae3fd6cd7b6324df10c3e0dd9381b353872af7d00d54f8889f12cfde9a9d1cb5eb0102b2c33f68e731c1546f38fe1d5a86, 512'h13b4f10be35d29df6da2f41486e5d99a7e55f8b095f8bae48b49c6dc69b123ca5baa15bdc29147023a19bfd6aa2e7aa4b848b6f4de5e6a308a5454c7bf82435e},
        '{768'h0c59569e12501d609f6d1a0432f9b2a622f833d1aaa20e87733db9070652cdac76f8c1b5adcaac5a51da78ef849b28941480ce0727fec6ee302b37c76710432b2ca7a096f2b36768d0020b69b39d1decbecac7929457c7e5f44c2b0ebfcac9f2, 512'h2c98b3a2cfd8fe71475d0983d2bce772afba63ac5cdc2dc09928bed1562a86d02ea39005b82e55070a5fc951ef29c14edf32493fede00fae9562b3eca6c9f032},
        '{768'h14b71d2602c3153738a0b38fc80f6e8b3dbe4444f5a906c4c0cdffce625c99414d4d85f90cfd648143f1f5dcd7eb3c83bb3c8f989325085fe02092d4a4af635a4560f1e03667a040a2885193e9cbe9842be64d264bdaf38295882d006f305d79, 512'h673b71401c92b2741a8e2c7c1b0cf61df7007e72fc369ed4eb1685472c7b144258c050f2f30d55f8b875ceb7805cbf16657c50a44d22aa7881d33c25d38f58a8},
        '{768'h155748c18950cbce663a9b525865b561903edd0892f4e9e0d38574c3fcc4114c333a9ff2e1ba968be8879ea70ea4bf95eece31d0fd0785c5812d005bad583971000f1453ecb872729c874d5f59502d43c2d22bf7156d192e195b433974bbf8fd, 512'h7ec833284b3774ce89098c4206c71c9ce69b876dce24b412472d250e0e82fd084d563de9351a5f330ab5532ad8333b15c5f85ecfe6b5d8e2114211f9da308a80},
        '{768'h5950e756222ce60e12fd7a65e9c6ad438eac73dd11434066d897c926c589bdb965e8c05fcc60be48849277e8b66fd92ec51fd69c87b2bf25d21c3cea887ae6a358ee438fe9470913f0a9acc51b7b0d72925ccd861e26e61d548dd963d271d4aa, 512'h7d949fc400fadee371deddc8d804a7e5087fd3e1b8a2d53a95e841fdc5d13992453b8b956a84d9560591e346c9b600d3c1ddbff585d853157a59fd1767110ae4},
        '{768'h16ecd6e94140de7b05873209d479e062944e0f1309d0edbb14e33ca621ae062165ffbc60468ab46d209a069da64f5ed78886d31b9c7ffd6cf7d62d80a3810a6915630b7b71f973137fb1141ff9c5a9cb4ca377912ba34f6e4396e9863435af7b, 512'h10a7b981363de48f4a28fd4ae96c2e702485c7c77c556014a9fc32dd609cefaa72533e761f60ad8784e1c9778c755ceb36aa16f7a29315b07ca488d24636e8ea},
        '{768'h78b3a109983b65705e59952859b3a56f1bcef2604046e14029cb558c5b9229fa3d797517d8ad8ce4d1a0803636f764d99474bf3817b4a7ce50d353197d4822620c2263e0d3d95ff95d003b4787a75843f7d69ff47212d9939ee2194e47a665e2, 512'h17ddf097624a1f5ef60216f13f06bc5772e52cc4cce126ebcd4f4779141e605e5514b94375549edf2c16080445bdb7495a07c72beb302281c168f326ee38c5b0},
        '{768'h7455ff17f4bb6cbe3f7d4cecbce13b6b8092cc0f6ddbb07016a9285c6f595a8f441388913239f541f18e6f54899ee64645ee0ed7f1966c4c361d289d05c79c840dab9353e1265d50a21f0b5eb4c1d6c04520ad9a4ca43c9f551fcd472b1d0cf0, 512'h37d0fb04a1cd688221732aaf282101640d3aecf5d8c65919686b469ce76a1f00158d70537ca46a25e3728748ef62beb41688214fd68c04a45e9e3cc7941c4f62},
        '{768'h471221d191aface80ca8e788527b66f08a7752693bb9048ea9a63887c7d3f2ff30d78d2eb628eccc956daa1e52c4efb43e769b0c79070d53ee5f10c7b8bbe5c23eeae667325cfcf5cd2c9f60ca4b73b2c79f416c527dd7f9012d44d9ea91160e, 512'h7d333e1422fcd5b54d25f4c61e3080c0a5fa75d3602b9f21fa7322335af35cc2571f161cdc708424f35ad3e916f922469a9cd0182491e7d7a8c60aee490a196c},
        '{768'h2755d861591765d436d3c0e7e19d90df006ab9efca258f45b802d632262d360021288982dc09d98065e9b2c4237b21e166a98f21ee1fe3e38eb1c99d7b5a83b345274c6c2ffeb908047bfac7b0cdff7b8ac5dc1010be72e55ab2829c3bce4cac, 512'h32d8bb6f8b3b9ae6560c054c75659b04e7791f94a0aadb1b28f0ddf64342380e07ebc14d815580f0cb204da6abe83c698b4201ae0ee13964fde57f5ae2fb5646},
        '{768'h55da8ef17a8ec4b54078799adee7f74f78682a32ea0a923e5f983f4fffa5751421adfd8843729ad90e161cd776bbb8aefe155d2ddca0b7696ac78f959667adc11a059f53cacf95eef76a35b5a20fa21d812b3502e012b50f13114533e2204afc, 512'h13b5c4df60a4d5501bfc42f6d7765aa698e799f8c30115844ff0772d289232dc151783bbdd14152b4b77a3da4f904efa6570bfc737e139800e30325bb82d6fcc},
        '{768'h3208e9a08cf0049064930741c01e82830290bc225b34bc7941ae603f2ee423df4272beaa5ca2a9631c4fef256df8c4323c3cf89d4be4f2ef069decbac7cf9e8d32addb662b1a1d203442d1fec9446e12ccfd242b014cf15a1f1da1232bd46beb, 512'h6007fcf63f18f737202ce5140e33fb2848e6c982c378de948b1869121f161956724a2fa7d0996ab5dcac0e4ebe94ede567890aee9d2b338b93b96d661e43844c},
        '{768'h13978703522098071a59ec2c0f91191dc030dbc8cdf4953e4d94ff8f137fa70b6ace5cec59d2a8ba43bc7e187a17ae861bb1a7b7f750aa1d3e49d3eb32212d0529b87e5a64be184ec0549ec5131d464f10c3dd8acfb8164432fb31e795834907, 512'h3791ddcf0d806ff4b50c463bb8b315e963d829d9a305232f328367a4ab7ab1861a20724114098fb7d162b106426d2e57a94127e831499972960a5e6aa983862c},
        '{768'h6b4f12b4f96e581a6030930f57b0741d0f3df47a106c9895f4edd696dddd551236f1dd923bfa5f9884570d866ab0692c9a0da3ff152d293103652cc1768ee34f379b166f6c27dcb7590280ca08b5e6ac2fdeb1580fed2be9c2300ce2f306b12f, 512'h0b420552171066a120a66c48b9ed4e2ba04e5bc3cd6cf8667b395ec221966558288661646a8b47a1933fffdbe2a592d315a783d01e6213dbf5d7af0d2eadc578},
        '{768'h0635b3174652cbf71bbec451e6597bec77daaa6100ec2564db97a130bbfc30864dd9673d16766a884ebb328af5ab996e7895440c7d2cb9ef8d7e9ff66b817b0b2b796a3797c5beda2a74533a9172ebc0d5d1ded5924a19d4822b6705f4688dcd, 512'h15cd04682a7f321248f3b8d10f4a23f84bd5e7d48e6560f6e73d978da8e9900c6685f6c92dbf8c648b3d9b40c20e9060bb661af0ff411d76b94ebcd4495227ee},
        '{768'h7e0488d0567b98387c76e28deb7b26e4bf69a395c06f698b521febdaa3365fdb68ae81256cc2f99699bd8ad6820df5cc0654fb6e6ddb79a75b859387315edd4d0882e6cc8b7fb60aa172de18c36238b3004038b25d113a77ba5578fba2f6fe73, 512'h445e265629c7d24745ad70e281683a3dffa743842d3e210349a990fa79b0afb21038c3b32368b4755062d7460f89cb8686334cca0c7787af2ae9aeafcc86f0bc},
        '{768'h443c20e491e8d9ac4160934702647a035dec5ad6000991622b7927414156d1d25653e01f4151cf0d07c75200d8831c4717b57d189e4a6358002cef7b54965c3766f41cf73569146412acc0485729724824d1be31607699751653be23727c3748, 512'h1603044efc9cf74475b666fda8a6511099182011ebb41a4665b0dfc31dd902d06e3be97d62664dfc6247a70c1cb3fd22693b873e4df02702150fa3177499f9de},
        '{768'h481797f38f5f021d829660c9b876a244d6d47adc7de95479f78837247539a58a188aea7cd81d7eb5d0f542a039beea36c31877ae376dceb5051fe8627047715731bfad0b093f59c3be95e3bb25554f9cf8ba0264f2eedd4a7921678742fe5a1a, 512'h0c92754475c7ef0b42489baedbea0a1d97f841972d4865eeed75f13696b0fadc323a7a5b8ea97aa9b08c2efbaed0ea10c1c21c60c4f3b96242845552229a5e08},
        '{768'h39d9d0d0ef67b01e34388cb63e9ce584909c975cf2de554d3bfbf3e6cb18b016046b8725e3dceca4991763123b15b172be0e977f383baa9d3521c6135f36b11447fda5259abbf0c44f5d30db1da782bcd1cd0ae044562ba552956e2dc33bb696, 512'h189f2ed7c734da9f84bacc7b49a29234d52d20bf283bf21bbacffdd3a018aee42bc92bfec1efe064b965d95dabb80f3423ca6ab4b1abbedd98692abaf61c6d10},
        '{768'h409f5ac100ab2e0a1d9e918af651167c4b6829de8517fee49e600c8e068808a669d9ee4de10cc743331df49b0bd2f14c43fd1c905289448a43b9223f6b0ab02e2b6f0d48eac16296057394c9788974a1b5a215f7c814042974bcc38f62e7e33d, 512'h6d1b4923f7e3b57db37d865181c3a04ec29b79fbd148b777300c8ea8ef4cee58739605487386b92216e9dd3de255d666157ccd73e9fb71dd177039c4e7174384},
        '{768'h59ea74df98145ed067b5ae06b527db48b2b12b13a796c2c6487a5f3b3295d25c5ab62bfb1d73693b6898bf0eb3fef3985849cf926d008960a001e06c488e787918549c616ab31ee8d9e4bae50217ab366b654e0554f34772dafe431118d0e73a, 512'h7b8ff41e4d405996244ef081a567a4b732a17a35c49b1023515b82b8e705f8b43c5be4425c3b606135b989b51586260511c6fccc972d1a274bc535861c16c5e4},
        '{768'h1695286cfe200915fa844abf3da7460bb6460b6fbf34855c6687b503a4ae61ec433ee8d07df09ede9be6d3616dd2c451e2cbebe29e63508aab6855111eeabc6f146fb0c64d23f524879fa8631c03adf1b28f75d26904f492462d40a1e0497b0b, 512'h66f5ebc1a34aacc4d3d453f90e546e42073fc0138d5605c4bf5c6f94eaf75ae055fe2df9af28021e2dadbb11bc3a99bd40aa213a20ab71b2d68625fddfe7582a},
        '{768'h39b590f59c5495fdba8194fa21ac15606e125584f552496c978ab1866b3ff7ba61e68f914941a9b8d2c38dfcc04d2cb91d948dbd0313bdbbd12fcad69311e61b48658958887943a79d96a22556cbf427baaa51838c599508567048753fa425c6, 512'h5fcd67dd92469da405b9e36afc87d59836fc8333b8603a2686a08acc4fa84f6610ef6d0412a284b32c4c9c7972d174113cb28e8b05bdcad4339458a05e89a60e},
        '{768'h3952d6b59dfe972819d3e1de57ac5724da0d9e7074a5a7af0bc36afd986a6e99632bd7e40f09340ccfd867f9007677f73693a1416e57acd7646bd516f9ea466965d2b96872a04777291c9dcb871ca1b1430322096ff17c9fccf92e8960379001, 512'h4101d1289d4c56bc927dd82daedb349a99467ac415cdfcddb4026d9e3933277025d5fa06bc3c6c2ee3fa2fa16a82d5788acc25f79531e9393f7daffac7d5ff16},
        '{768'h28a7e7a714ccbed4103aed8aee338ee46bed1c392ec341ed5d4f42389bcde1537d6b485025a0a4b1b21cdfaa5235dc01061e860978bbde7d328392df1fd9edf277db6290fa15b0df33f72b0cacf5410738092c6e629354b70323ed9c0db92d00, 512'h2035ca13bd041d2687026e17970e02ff096f13dc299993b89ca72e97edab3a4c6fe6f0c91c81c2b7838a450826ad1b4649d9b9c8d2f9ea121647137195d1f638},
        '{768'h026cf3fb57dcc43f3e077875d43ce247e4250ef2dac1295ecce76da942485a425811cabb8e07327edaca6ff07f10065b60463c5af7e9d9157d5ee5c527ab7baa69157358a10ff24dc7d8b4404a849559bac8b2db78730d71394ac683ea9ba422, 512'h609485e156e71064bede10e9d44fa2e68c15e38f8fad26e75ef0a5496051e29c3b05a086e8635e342fdc3b53353950fd38052e6368a59c27557ddd15f28e47a6},
        '{768'h404431b06102091b85058a3b38938c756206b4807c60926a0daf21686b44e94662b6ce903dffe3ea6c7e0f98b303386099149110fd877c7f55e85b6d41dc9992064a186054ac7c6745a2d64409f03bf4a3083476f739199f8fa56d2e89ce7b47, 512'h7a7b39ce23afed51deceff10d28b3ebe382b736a5cd10377ddbe2373de42345214692a0f6a1160557496dbfeca6414db8e0ee02c0f883a3c5e1793d139d34fbe},
        '{768'h4525dbf50acae6b29d1b0868164c2f7ba27537e808ef602e57c1e4c0c652662a3cb0778705d67921d21eda754ea7930eac2d4dcd1e1bbcceadd354b523d5ca2c0a49ede3939c8968cf9517353f8d5e9e58dd786da810780472ca50d67fb3cf8e, 512'h06c4379cf1aa95f6df6e8f23ed328ec05c28e367f0202943622935b60135e4b207ee67c84af6e7246d0d5b5c9cf87343fb699998ef9d81e114cab8c3903ee824},
        '{768'h53a4708c44b5d39feb1ab801b50275d1df03568f99793ede7aa15f99cf8f7a9c63c8717cee0b42d645ec85d5aa35d4b0b851a7dc7f9d976493592e3158ee0afa3dded8451be0c429a87e4a897722333d943ecedefef47c7f2c3f78c3779484d5, 512'h71d42ba6be7f1ec7955c1047ed0f1ed84056aef26a4384cf04be267f2034667e7c2a0cc36367d90baa346881ce02288587d51e9b96d547f56c0d443ce2fe34e8},
        '{768'h5ac6a2900bdb28a75ff2f7758c13ddb2d1dc9f02c89686e75b05e49a05be8dd50dc0166a072b31636d3c4a40b6264afff16038e1220159242de6e6095574645a714cd7a12f950633142799d7479cafa4e77fca4abc6542b87ccba17fd68d401c, 512'h30ca9efc302aa4ee3eaf7e53d16dbe9730db22a5cefcfb6a5f4f5c312474c1327a0bd2040e00381bb51d25accbf9cec950c185525801359e243b3980805e86fc},
        '{768'h44bbbfb4ec25bb94d6d1490d8a80ee0f7e1c75850e6cc4760504b090b55d54f667a3533d30ecb3b1fd12f3b6a8ab99d19b51e73c1a48d3a0d18acc8ccd9b41d7361d028b8348da06ab8ff6772469181107c0ba613c95b2d403ae1590f2c43812, 512'h7399055e28b53aeb60a318f01b193421f9468ebe4aa674ba9ef90a1b1ff631f4051080a778808cb463a0b2ab1f2af50f59609c228582ac782dcf0d82f54fbabc},
        '{768'h2e9ef7c66bbad242fcbf54e0f47c0c4fc0fe91d634bc12ebade3df70f9a425a465aafb18ea8b7990f593d4ff57bd84cac28130bb3841e77b8a8c1e28d6631d5d7ce1fcfd8d62ad492dd3a5a7256bceacf6570c46d69330aa27e85d84afe93744, 512'h107bcb128e476ff6491642bc9b1bbf23498fd8bdb91411fee7bd75f0c86af98052af7005c6bc4517b3f1bc1d32b3a6d36360ac721fcbba8697327a3e91f56fb2},
        '{768'h4f967636bd1c38caa5536f8412310ab3e5eb9604ba350b9e9f8ba8f666f143ac6ec194400658cebeec7675f060a49d8ad584172e7d2aac59cb61a2a0b517f0563708e56539d6f4a11d3804abcf608fa58f24e574213e459b0f51da0d19a18173, 512'h4df86c2f3e5814e1b164d0b23799cafd080b58bfaac490fa1f82ab3f80dfb15a06e456b8d81485905dfe4ff74211d2381f39f12685ada6ff5cfa94023fd4d332},
        '{768'h7fe3a4dd643c311b814972c8823e1fd2a4f71ca9eec80ef32747b3bddc4e22395c3c09c2f96295b70221839f44ecb017afa5ab30c8f5ec8af15c0792cf5f1572716843f932eb3f90bd9cde9d0123b57fd4c2c3fb73d1978f839df5dfadcfc895, 512'h2acd7ebee95d4b386ec95c8ec12b520bc26d74228ce6b7a5ba391e9219bb4ff82b79542293bdff976f4acb4f76922e9a68411cb07ee2be2305268b3f866b1dae},
        '{768'h7ce500ace8662ecd092b3b952849e69ac2070a392c23505691f377cfecca55fa666965a4147d6a00fcfafb90c835e295749cdc4b1f6436039e84c8aaaf469a174d8e9459bf76f97916f0e0db76a031f424a92f8a07a9af00ab504c55327fee77, 512'h37cc2f090de0fc86b1b8087ee2b02c575cd0b181351cee661daf363bcde1aa404fbbd68ff94459be572ea26108f4977a0bdee8439b27508dbdb12a88f1d162f6},
        '{768'h4c912069ce4a1013c34d8f52b6b29c729b24a7b00a005013d912c0be05638caa38b1477e4679ba557262b5ca24c3d0e85344ee98097969d566c9fee1557721d0116b27c675836f178a4f7e3ceca4b37bc538209c1aaa3c26447e6135b97502f0, 512'h3f3d63cada3ebd6f852df16d9aa9006a3524209570842d6993325a617237de14514010c6416b3eda57f3a5627bb5751a005f5421b4f0b13bb6e9b6f584a04392},
        '{768'h1ee698caa0929089ff22b257c555fe9cb6eb77c14dfd0e697c391c4247772cee44f647cfd1a26f6ad4ec376b71999eab0dddfdbe0b444c2a8c1599c2b517ebd7187604765bfb81395293bc16d866cff25d7cf3e155b04f940a90c63cfb214c03, 512'h1a6d2c01f4ecc2be0178c744aed6aefb73feb7c457a62db48f111499d8b2f2861da9859b83d397f185864edd38fcc9509cd3f0e4766275809e592a93b53ca6fa},
        '{768'h51d2955dfb55875314a2a22b355784dc1d1dc7dd5c1b9910a39f5f6651a6c0d34ec8994d38f6f0d6ede8b29f0fe42dcdb1f05deea76992d1d8b4d631ca06331c536c35068efe5d28da091ebb8484dc749709fec4fd7b69b00c04ef3b9e6d9029, 512'h79729ce758e206caa8555f0a35086d5e4cd6f952e21d25fae6e82fd8d2185af84e47133dcb65727243a481eebe28538a90684f834ff7bc9399a5123d3ab68940},
        '{768'h1ef2f9492ce5fa91925a7ff3751a82fc5931eb43033027e91c02581d29d114a957e3c219add3590afbb53055a9f0771cf5370b52df2bb6a1f49f7238540ce3de1e4fb6b2ef6ae9ff4373679b91eb01525c34a7bfe2e31a7c49425f85481e939a, 512'h3e000cbf7082e1efd709c2654505503620c950022ad882b9ff7f9cd95b47006a680de54c51d1445aa8c990fabce483ec09a519ce0fa6b5b828ab6b40407d2260},
        '{768'h3f2b7ba55d51ac9b13b0d61b87788e40c13c564b803d9f0e1b9356eb47df19d51e9d1c57b889c4543e502c15f5e63a98596a34a593596f9c313e355670b593df7e5df472a4a46dc682011e609901898d5ad0e352e5b3241453221a909bb2dde5, 512'h4ebd00b2cfe4596697f3fac1e127479b59a202de1265a64d90f7d7c6512c6572483d11e4f676ccd936d9fffa72633910a2df45a6a16b842eb286b710d9cdb7a6},
        '{768'h02180ca3fd3ce8dd1e48fa4a626c4a2d95acb3e175a27ca45132d081d5efe80967f9974681de5978d570661a2d09abab3bb12ebe4f67be964e5a19d53d4265594c329d98bce81c3c4d2c2571f1332b06e85d80d0b292cce89772b9c3da441cf7, 512'h27eced91f2c72590bc833491c026bd0e9ad9961470c2ef91f8ce82b0159317fe76b359307b29b6a5f30534ebdc75e7f8d2ab88b44ee6fb81915527e4288c386e},
        '{768'h5a24b7b36f8c7f75938d0552010ef24c498a420b35d579baa0261ce8d764cbed6d47dd24aca3799e644c79211b330808a0ba4c6dcc55dcc8de9bae4c1cd2bed0534fe5524ce16240ea0cbb59157c4925b01b46a1a2845ba5742dc8c1328fe873, 512'h3bea8dc7bae2e44869fcb68dd577f310db59196c65270274c220be19a74417ce7773504f5410fb663f84fb4cc7ca82b04a6a4fcc166d6551bac2bf23dee82af2},
        '{768'h401d8370f91f9d4c3372a4434e8c2a532f0d0a6b14b7b20aac6ae60260cfd1df2a96e206e16dd6b4bc50f27f261e44cbb5cfea7a7cc47f7b6b6f098d1183b31866b88f8991d30418778254ba54993af42088d93cf5eb6d59aebaf1ec5c5a0cb5, 512'h0083b42b00a925672512e382e485694323e22b64374cba19ac7b571c2471cf6c58adce9a3060b85843b3f37de368e64327741dbf0164145261215fa42c06faca},
        '{768'h5e1ad46385a8d1f295e9de9ce4b91c032f1ed890894a710fb7d66fb6b6cfa49d33369f66eca6e6cd3d213a4a64389ee77850323f2b4e08da34b41ae694929d1b1fde9ea472bd0ae18b695d52fca6bf5335c9e4eece9fa8461613ce29a5e67c09, 512'h74cf297aefa015731a2ecf71474603cc8b0553903c98b715cce7fec130a0be700350798b348f3b228aa1ea874fc1d12eb9c7b9ba046dce85bbb2c9c732ced93e},
        '{768'h4cd75803a8c8e4d040ce399897982b6d79880173009dc046320a23b8b7118274221e02a25a04eb944cbd4354ed3907dd48326bf6188e3089ffbe14f614966a224631d12526183cc8552d3cc756bee79a7af44fafd303d0a33e3ea9d685c6d920, 512'h42f1da41cb7ff1ca4b4d76153c9e4f16a05ea2f26aeee123ecbdc150f68a4708488db64b7347202d69787ceee051bef0764056f24fda2be41e09820780aca3e0},
        '{768'h221e736b6112cfe68625008d4e46514207680dcfc7687b2be7179d817a0ed98a401262d9f8bee00ff0f7b0898a6330ead2a754df2591f575a8130401834899e5123105909b77519c89e17cf9450599f1fb91ec7fa6ae1e27abb0b6d552b85ed6, 512'h370db4af0ac2e305c5fb4cd12c095a99af9b96cc25822a31d3cbea20927c48bc354acf255f9e41100e4e03012424b9572ab84a9cfc55bb0bc7a44279f41725ec},
        '{768'h64697f07eaec94439fd15583f03879d062ee3cbc3cf3d77a14ff6af7862b176517909ff2054e9fa9a7a6a065ef4f46e16fbc222c3d565dcbba376a598732d95c6234303d65f99ee231789f1692f584c68481acbe4eb4f5a9ddb49595b09aa381, 512'h0043cd4d1c66bae50fd4730256742ff2055fa65af5670d5432b7bebea1d5160065f8ddc4b90447f70d23d467195d29d1835944377c591c9be7ee81b6206ebb9e},
        '{768'h180778e96094727a08a798f8fedcf57ee9712d1d7fad5e2886ad35e7e42873ae32758e5b9b28259b9d21b2e5a7f0ffd396529d6f977dc8356a274a6cb6c9a9c0151117df16b77b5a0a5656e4f8215de8ea65f50d7ec4c3d6f6990471063467fa, 512'h1d98ffb1e93a738b49e728b86ce906d18e693d3ac8ce3e21536f04b84764a99647f036c55cb5b3d350e16f4a3ffd314f01f040b6c1ef23b824123b033706857a},
        '{768'h79c1a19c3c55e1406c2638631ebab1fc1d26aa3478d6d230ef8da4f0b0593bb634eddb3a7cb46034c789e28d6936eda531413860096867fcb7dc1d99c54ddb6c7d44e326c7c290b15f1875cebb634da2dee973d0aa43f18f5049869309494435, 512'h74d7cb9a535661c605d31ad24e28da814621e645e0a8a72614fdd10212e724843375dbdcaf371d6a34dd580aba668e5ccbb3fde3888f14d2d8cfb05a26edce20},
        '{768'h2c2cc2cbf320f66313d1237a7e71d8d64fe06a38ad8381b2e5413b8598893174789c738b9c747ad4ef15af1a489feaf20fa0fc61f4fbd9dbae734082be09f6b130cfb2605907d9aa485aa2535c59e0cf110dc101188585d7fa97fca244788cfa, 512'h0e5fbc51ee8ec9517aaadf09e0c7689a7b8ba5df9ae4c239dca704e35509c9627e9fb6e9c63657b7d544cfba45df91bfe031f75dcf75cb2e802e0372ec05eca8},
        '{768'h14b92435b47156e98a74608aa2300dd5abf6098a54da7596fb05ef78f2d14d737ba523b8f4d3133a5010df67f985b083fdd9c44f4f40754bae89e016f4fa635731a6e5443023a606cc3171a56c14dec4bd1b3c55fb4ba30467175a27deefd86d, 512'h770ff9bd42443ce9168f3e776a87721ae7973b76d0ce28a9908ce56cc92dd1d8786bdddea47d605757d80bf0264e2935baf3c20a39b79494c59d0e9d1206c812},
        '{768'h487cd57ca9aef5147cd50e72708ac2776bfff98110f428dde1554071f8ff8a475c3601124f53c4962098b79b4d8c28ffc17362bc20a139afe43c1eb83754b93915b71b737a63f7879863071ba84ba6ba7255c53757d66b9db9123cf7d214cc09, 512'h063b1486dad500d27c7c75d68cb0ff340690c06bfc2074c30e9ebb3d4d2b426249f52ac0a1c23a3cfd79d26ed7f44433e0e9026496afc47afa0845bd681b598e},
        '{768'h27cf7e36c9f3cebb0fe1a79c97ab627a1f51c63240131c5e2030b49cb156f48b6bba1d034785a99c39222855b200eec03f73e80cb824810c796c272c79c4776d7b7a98f609aa88a8d1517373e32695fc17a65bdd245e6680f68a9f3ca4d40aef, 512'h142635c7bc0ea3f2a3bf5bde1dbda9c3bce0c5763182b9af7cdfb2a2fab7d0ba136b406f8bb7f03c5c9f97101aa2667085b0fbf006a108d4462ef335d3b2eabc},
        '{768'h16438c365f0da961a06ed61ea1696885c71167aa88d2a5a071a7f84e3e669160177a9b9d37b31162559b342074c12aa5697ced420f970fae5863747e63f82bbe3a3f821dec65d2e175ffa90d24d3f49125551c4abf962952cf3928bb158debba, 512'h3920b1a600baae56b8a1113270d62f607f369c3973d86726a4a26e23861bef84731370217dad26b120e741408ed6a302e9c77d8cfe15381a55cbdaf8e971be5e},
        '{768'h392666da6c5e203eb64944cf44a1eb02187b67f8751a6e381862ba7bb6ec70b77fa0367f3794e5df12ae9daf02e309a7bd13d9441ce88b0320e2bb2decc4aa6c22058c0570967fb6a441e287d5820d3cfb39f04c08278a9e7f26f684edf7a293, 512'h6aa986cdb54e4a72b5236c94af8c0da1d4b344686d9fe89b280f7c090d1f0fa242a86d55826ca92f760d105d30eb24a9ee6b37c9ec02648b73a8dea697d9784e},
        '{768'h322649aa0d8b746f98b737521ae1d453e3b5c9e0de0e9913b42fbe9804ebf93f25838f6480b077c7aabaa474a15ad3ad010f06a4b4c72f1c28756ceab7c81ff86ba5f4078aae514090f9e6be4059fd8d2092abc0bfbc10b2968c6a28fc1b0892, 512'h1a4e060a44e1500148d8ffa6347be08e4a0b8567817fa8c7909eede2191121d41ef0682acaa63267013ce3bc5cf5a3797dabb5c1da2fb3a98f32eca81edb759c},
        '{768'h3a8237f77a07a8cac94c67a5c5f3d24f8b22ac0edd228e2d742dbc5f9dba6d1961854ce2f40ef201303e752f35e3e5465ac6ec95f1c378a71d1124c5a64fd67f4e97654946f5c41ec00e3eaaf23ad01b7dc171e11ad17c5c32496319f28dfbd7, 512'h5905d49114817151348529651c252f8706ebcbc9b8b323db589ff108d39cc8fc606785e84355642e7a6bde38aac03bffb972c47e4c3addd7f703ec4def56ca78},
        '{768'h35f1f50b7ae1178fb7c3cc64b35306097f2c5246cabfe7284e88c2589e39e74220ed6686aeecd91198d6544908d1b27492906968f85170045c8aa0d16f7c8e376264a687907bd4957a6cb5d87c340de4c0af5521f4369296fb6a95c475de366a, 512'h69fc7e96021f5973bf618d21cba633d01c5e2f37fddb01434eedf5e967055ada3d9c7f47f7f7e08044e604fb9ab070eb30947d58cde0818f091bf57895e23b96},
        '{768'h2469f031a65ac7199d9bf1be4fe6359c6b642a05a5a76d307857f38fa28b7a187e6e634cb275cc698e635143c56fabadf3ba872aa68ea9201b4c79ff10a9c8c55bba6a5d3937c390d1b0906377bb64f54f7880fa4ad4fbde92b7922ea367b151, 512'h594ccb89af4e5abba8d705db9b610b4005d22b847f0b1f62c0c57ea4ea6659a8067dcdf371647e51aa32b5d3e4dae0f5514b9562ce9627dbfceb2885e9d9299a},
        '{768'h7a18a1d405f9acd504457244347604cac35061cb3cc7943d686be04f52c3381a5e86e9c37b13bea5fd319573c985cf9201c4d15d86917a264f414b9dc25319bf64977acec0bb2fd5e97eb09fb1cf9d8ec13fb77ab4e81d700c4148c0d9d55414, 512'h592f94413348edac7f6c6b45557729fa3f01469549a889470ddefe57ef9784fc0c709546da523268077df9d9f7b98129fb5f565089f6b7bbf101c3682d80885c},
        '{768'h2ae95e6ed5ad3f0b973871b9fd52312f769c035162d5a0e76615d3d80fb5847d21ce97e22c1a1aafc2b1d1668fc497c9e5c19e715f9a88e95310859a8e4a032505303cba89b12eecbe22953cdab3bc62980e959b714e0dc6b43c31fbe81d5d3e, 512'h6d32fddb1f69635e554bf760648996e168125f7cea2e0202ae6e18736d818db24cdaae3f971156259e659db57212c5328f51c1dbc085ef2a2fb3fb02a831502c},
        '{768'h20051be45f046198f4fd1c59d8e7411afaa89cfae528bcb71737d786076e20f6697cdac7e2611a680919c8318abb8f012c28adb3119317fed8960a90fedf0cfc38bbb5aed27af310d30963aa21258b0136aa18cc7c38d1cfaad11d40cfb25b4c, 512'h4d1d7210a62f9a867e4c07f3901b353f9580fe730381126b521ea9b26435498458210145cfff1a175e9aa26d880b2f1d3240541450e20de44adb0fe99e2b16aa}
    };
endpackage
